interface WRAPPER_IF(clk);
    input            clk;
    //Module Signals
    logic   MOSI, SS_n, rst_n;
    logic   MISO;
    logic   MISO_ref;
endinterface